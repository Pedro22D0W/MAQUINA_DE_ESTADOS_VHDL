LIBRARY ieee ;
USE ieee.std_logic_1164.all ;


PACKAGE CPU_package IS

COMPONENT fulladd

PORT ( Cin, x, y

 : IN STD_LOGIC ;
s, Cout : OUT STD_LOGIC ) ;

END COMPONENT ;

COMPONENT ADD_SUB

PORT ( 
X, Y : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
Cout : OUT STD_LOGIC 
 ) ;

END COMPONENT ;

COMPONENT REGISTRADOR

PORT ( D : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
Reset, Clock : IN STD_LOGIC ;
Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) ) ;

END COMPONENT ;


END CPU_package ;
