LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
ENTITY BUFF IS

PORT ( REG_DATA : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
Rout: IN STD_LOGIC ;
OUT_DATA : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) ) ;
END BUFF ;

ARCHITECTURE logica OF BUFF IS

BEGIN

 OUT_DATA <= REG_DATA WHEN Rout = '1'ELSE(OTHERS => 'Z');
 
END logica;