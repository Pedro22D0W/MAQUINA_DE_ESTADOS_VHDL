LIBRARY ieee ;
USE ieee.std_logic_1164.all ;


PACKAGE CPU_package IS

COMPONENT fulladd

PORT ( Cin, x, y

 : IN STD_LOGIC ;
s, Cout : OUT STD_LOGIC ) ;

END COMPONENT ;

COMPONENT ADD_SUB

PORT ( 
X, Y : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
Cout : OUT STD_LOGIC 
 ) ;

END COMPONENT ;

COMPONENT REGISTRADOR

PORT ( D : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
Reset, Clock, R1in,R1out : IN STD_LOGIC ;
Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) ) ;

END COMPONENT ;

COMPONENT CENTRO_DE_CONTROLE

    PORT(
        Clock,Reset : IN std_logic;
		  FUNC : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        R1i,R2i,R3i,Ai,Gi,R1o,R2o,R3o,Ao,Go : OUT STD_LOGIC
    );
	 
END COMPONENT;

COMPONENT BUFF 

PORT ( REG_DATA : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
Rout: IN STD_LOGIC ;
OUT_DATA : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) ) ;

END COMPONENT ;


END CPU_package ;
